library verilog;
use verilog.vl_types.all;
entity REG0_2_vlg_vec_tst is
end REG0_2_vlg_vec_tst;
