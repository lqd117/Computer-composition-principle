library verilog;
use verilog.vl_types.all;
entity uI_C_vlg_vec_tst is
end uI_C_vlg_vec_tst;
