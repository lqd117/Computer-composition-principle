library verilog;
use verilog.vl_types.all;
entity uP_ROM_test_vlg_vec_tst is
end uP_ROM_test_vlg_vec_tst;
