library verilog;
use verilog.vl_types.all;
entity uPC_vlg_vec_tst is
end uPC_vlg_vec_tst;
