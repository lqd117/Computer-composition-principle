library verilog;
use verilog.vl_types.all;
entity decoder_B_vlg_vec_tst is
end decoder_B_vlg_vec_tst;
