library verilog;
use verilog.vl_types.all;
entity cpu_8bit_vlg_vec_tst is
end cpu_8bit_vlg_vec_tst;
