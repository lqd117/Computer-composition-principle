library verilog;
use verilog.vl_types.all;
entity REGS_MD_vlg_vec_tst is
end REGS_MD_vlg_vec_tst;
