library verilog;
use verilog.vl_types.all;
entity decoder_C_vlg_vec_tst is
end decoder_C_vlg_vec_tst;
