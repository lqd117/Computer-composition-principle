library verilog;
use verilog.vl_types.all;
entity Simple_Circuit2_vlg_vec_tst is
end Simple_Circuit2_vlg_vec_tst;
