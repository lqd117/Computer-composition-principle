library verilog;
use verilog.vl_types.all;
entity lpm_latch0_vlg_vec_tst is
end lpm_latch0_vlg_vec_tst;
