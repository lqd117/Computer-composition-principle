library verilog;
use verilog.vl_types.all;
entity Lab3_1_vlg_check_tst is
    port(
        F               : in     vl_logic_vector(0 to 2);
        sampler_rx      : in     vl_logic
    );
end Lab3_1_vlg_check_tst;
