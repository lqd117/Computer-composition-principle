library verilog;
use verilog.vl_types.all;
entity up_ROM_test_vlg_vec_tst is
end up_ROM_test_vlg_vec_tst;
