library verilog;
use verilog.vl_types.all;
entity CNT8B_vlg_vec_tst is
end CNT8B_vlg_vec_tst;
