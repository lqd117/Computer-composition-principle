library verilog;
use verilog.vl_types.all;
entity Simple_Circuit_vlg_vec_tst is
end Simple_Circuit_vlg_vec_tst;
