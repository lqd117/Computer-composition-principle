library verilog;
use verilog.vl_types.all;
entity cpu_8bit_vlg_check_tst is
    port(
        ALU             : in     vl_logic_vector(7 downto 0);
        ALU_B           : in     vl_logic;
        AR              : in     vl_logic_vector(7 downto 0);
        \BUS\           : in     vl_logic_vector(7 downto 0);
        DOUT            : in     vl_logic_vector(7 downto 0);
        DOUT_B          : in     vl_logic;
        DR1             : in     vl_logic_vector(7 downto 0);
        DR2             : in     vl_logic_vector(7 downto 0);
        FC              : in     vl_logic;
        FZ              : in     vl_logic;
        IR              : in     vl_logic_vector(7 downto 0);
        LDAR            : in     vl_logic;
        LDDR1           : in     vl_logic;
        LDDR2           : in     vl_logic;
        LDIR            : in     vl_logic;
        LDPC            : in     vl_logic;
        LDR0            : in     vl_logic;
        LDR1            : in     vl_logic;
        LDR2            : in     vl_logic;
        LDRI            : in     vl_logic;
        LOAD            : in     vl_logic;
        M               : in     vl_logic_vector(24 downto 1);
        PC              : in     vl_logic_vector(7 downto 0);
        PC_B            : in     vl_logic;
        R0              : in     vl_logic_vector(7 downto 0);
        R0_B            : in     vl_logic;
        R1              : in     vl_logic_vector(7 downto 0);
        R1_B            : in     vl_logic;
        R2              : in     vl_logic_vector(7 downto 0);
        R2_B            : in     vl_logic;
        RAM             : in     vl_logic_vector(7 downto 0);
        RAM_B           : in     vl_logic;
        RD_B            : in     vl_logic;
        RJ_B            : in     vl_logic;
        RS_B            : in     vl_logic;
        SE              : in     vl_logic_vector(6 downto 1);
        SFT_B           : in     vl_logic;
        SW_B            : in     vl_logic;
        T1              : in     vl_logic;
        T2              : in     vl_logic;
        T3              : in     vl_logic;
        T4              : in     vl_logic;
        uA              : in     vl_logic_vector(5 downto 0);
        sampler_rx      : in     vl_logic
    );
end cpu_8bit_vlg_check_tst;
