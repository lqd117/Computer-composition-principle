library verilog;
use verilog.vl_types.all;
entity testbench_2_bit_multiplexer is
end testbench_2_bit_multiplexer;
