library verilog;
use verilog.vl_types.all;
entity Lab3_1 is
    port(
        F               : out    vl_logic_vector(0 to 2);
        A               : in     vl_logic_vector(0 to 3)
    );
end Lab3_1;
