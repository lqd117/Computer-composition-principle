library verilog;
use verilog.vl_types.all;
entity decoder_A_vlg_vec_tst is
end decoder_A_vlg_vec_tst;
