library verilog;
use verilog.vl_types.all;
entity DFF_test_vlg_vec_tst is
end DFF_test_vlg_vec_tst;
