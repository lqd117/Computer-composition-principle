library verilog;
use verilog.vl_types.all;
entity STEP_vlg_vec_tst is
end STEP_vlg_vec_tst;
